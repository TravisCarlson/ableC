grammar edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax;

exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:use;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:sqliteOn;

