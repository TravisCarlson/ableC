grammar edu:umn:cs:melt:exts:ableC:sqlite;

exports edu:umn:cs:melt:exts:ableC:sqlite:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:use;
exports edu:umn:cs:melt:exts:ableC:sqlite:concretesyntax:sqliteOn;

