grammar edu:umn:cs:melt:exts:ableC:yacc;

exports edu:umn:cs:melt:exts:ableC:yacc:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:yacc:concretesyntax;

